-- making a new file lol
