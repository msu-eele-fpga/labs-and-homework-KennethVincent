-- start of the vhdl file
