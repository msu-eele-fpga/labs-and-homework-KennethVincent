-- start of the fsm of the led pattern maker for lab 4
