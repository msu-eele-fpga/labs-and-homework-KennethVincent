entity aysnc_conditioner is
	port (
		clk : in std_ulogic;
		rst : in std_ulogic;
		aysnc : in std_ulogic;
		sync : out std_ulogic
	);
end entity aysnc_conditioner;
