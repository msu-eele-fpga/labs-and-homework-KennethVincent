-- start to the tb
