-- start of test bench

