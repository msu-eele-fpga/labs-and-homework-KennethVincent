-- package for hw4
