--start of testbench
